
class CoreDriveStimulus ;

rand bit RSTn ;

rand bit [31:0] CoreReq ;
rand bit [31:0] Addr0 ;
rand bit [31:0] Addr1 ;
rand bit [31:0] Addr2 ;
rand bit [31:0] Addr3 ;
rand bit [31:0] Addr4 ;
rand bit [31:0] Addr5 ;
rand bit [31:0] Addr6 ;
rand bit [31:0] Addr7 ;
rand bit [31:0] Addr8 ;
rand bit [31:0] Addr9 ;
rand bit [31:0] Addr10 ;
rand bit [31:0] Addr11 ;
rand bit [31:0] Addr12 ;
rand bit [31:0] Addr13 ;
rand bit [31:0] Addr14 ;
rand bit [31:0] Addr15 ;
rand bit [31:0] Addr16 ;
rand bit [31:0] Addr17 ;
rand bit [31:0] Addr18 ;
rand bit [31:0] Addr19 ;
rand bit [31:0] Addr20 ;
rand bit [31:0] Addr21 ;
rand bit [31:0] Addr22 ;
rand bit [31:0] Addr23 ;
rand bit [31:0] Addr24 ;
rand bit [31:0] Addr25 ;
rand bit [31:0] Addr26 ;
rand bit [31:0] Addr27 ;
rand bit [31:0] Addr28 ;
rand bit [31:0] Addr29 ;
rand bit [31:0] Addr30 ;
rand bit [31:0] Addr31 ;

endclass
