interface Core_Interface ( input CLK );

  logic RSTn ;

  logic Core0_Req  ;
  logic Core1_Req  ;
  logic Core2_Req  ;
  logic Core3_Req  ;
  logic Core4_Req  ;
  logic Core5_Req  ;
  logic Core6_Req  ;
  logic Core7_Req  ;
  logic Core8_Req  ;
  logic Core9_Req  ;
  logic Core10_Req ;
  logic Core11_Req ;
  logic Core12_Req ;
  logic Core13_Req ;
  logic Core14_Req ;
  logic Core15_Req ;
  logic Core16_Req ;
  logic Core17_Req ;
  logic Core18_Req ;
  logic Core19_Req ;
  logic Core20_Req ;
  logic Core21_Req ;
  logic Core22_Req ;
  logic Core23_Req ;
  logic Core24_Req ;
  logic Core25_Req ;
  logic Core26_Req ;
  logic Core27_Req ;
  logic Core28_Req ;
  logic Core29_Req ;
  logic Core30_Req ;
  logic Core31_Req ;

  logic [31:0] Core0_Addr  ;
  logic [31:0] Core1_Addr  ;
  logic [31:0] Core2_Addr  ;
  logic [31:0] Core3_Addr  ;
  logic [31:0] Core4_Addr  ;
  logic [31:0] Core5_Addr  ;
  logic [31:0] Core6_Addr  ;
  logic [31:0] Core7_Addr  ;
  logic [31:0] Core8_Addr  ;
  logic [31:0] Core9_Addr  ;
  logic [31:0] Core10_Addr ;
  logic [31:0] Core11_Addr ;
  logic [31:0] Core12_Addr ;
  logic [31:0] Core13_Addr ;
  logic [31:0] Core14_Addr ;
  logic [31:0] Core15_Addr ;
  logic [31:0] Core16_Addr ;
  logic [31:0] Core17_Addr ;
  logic [31:0] Core18_Addr ;
  logic [31:0] Core19_Addr ;
  logic [31:0] Core20_Addr ;
  logic [31:0] Core21_Addr ;
  logic [31:0] Core22_Addr ;
  logic [31:0] Core23_Addr ;
  logic [31:0] Core24_Addr ;
  logic [31:0] Core25_Addr ;
  logic [31:0] Core26_Addr ;
  logic [31:0] Core27_Addr ;
  logic [31:0] Core28_Addr ;
  logic [31:0] Core29_Addr ;
  logic [31:0] Core30_Addr ;
  logic [31:0] Core31_Addr ;

  logic [31:0] Core0_Data  ;
  logic [31:0] Core1_Data  ;
  logic [31:0] Core2_Data  ;
  logic [31:0] Core3_Data  ;
  logic [31:0] Core4_Data  ;
  logic [31:0] Core5_Data  ;
  logic [31:0] Core6_Data  ;
  logic [31:0] Core7_Data  ;
  logic [31:0] Core8_Data  ;
  logic [31:0] Core9_Data  ;
  logic [31:0] Core10_Data ;
  logic [31:0] Core11_Data ;
  logic [31:0] Core12_Data ;
  logic [31:0] Core13_Data ;
  logic [31:0] Core14_Data ;
  logic [31:0] Core15_Data ;
  logic [31:0] Core16_Data ;
  logic [31:0] Core17_Data ;
  logic [31:0] Core18_Data ;
  logic [31:0] Core19_Data ;
  logic [31:0] Core20_Data ;
  logic [31:0] Core21_Data ;
  logic [31:0] Core22_Data ;
  logic [31:0] Core23_Data ;
  logic [31:0] Core24_Data ;
  logic [31:0] Core25_Data ;
  logic [31:0] Core26_Data ;
  logic [31:0] Core27_Data ;
  logic [31:0] Core28_Data ;
  logic [31:0] Core29_Data ;
  logic [31:0] Core30_Data ;
  logic [31:0] Core31_Data ;


  logic Core0_Ack  ;
  logic Core1_Ack  ;
  logic Core2_Ack  ;
  logic Core3_Ack  ;
  logic Core4_Ack  ;
  logic Core5_Ack  ;
  logic Core6_Ack  ;
  logic Core7_Ack  ;
  logic Core8_Ack  ;
  logic Core9_Ack  ;
  logic Core10_Ack ;
  logic Core11_Ack ;
  logic Core12_Ack ;
  logic Core13_Ack ;
  logic Core14_Ack ;
  logic Core15_Ack ;
  logic Core16_Ack ;
  logic Core17_Ack ;
  logic Core18_Ack ;
  logic Core19_Ack ;
  logic Core20_Ack ;
  logic Core21_Ack ;
  logic Core22_Ack ;
  logic Core23_Ack ;
  logic Core24_Ack ;
  logic Core25_Ack ;
  logic Core26_Ack ;
  logic Core27_Ack ;
  logic Core28_Ack ;
  logic Core29_Ack ;
  logic Core30_Ack ;
  logic Core31_Ack ;

       clocking  core_intf_pos@(posedge CLK);

	      default input #2ns output #1ns ;

              output RSTn ;
                         
              output Core0_Req ;
              output Core1_Req ;
              output Core2_Req ;
              output Core3_Req ;
              output Core4_Req ;
              output Core5_Req ;
              output Core6_Req ;
              output Core7_Req ;
              output Core8_Req ;
              output Core9_Req ;
              output Core10_Req ; 
              output Core11_Req ; 
              output Core12_Req ; 
              output Core13_Req ; 
              output Core14_Req ; 
              output Core15_Req ; 
              output Core16_Req ; 
              output Core17_Req ; 
              output Core18_Req ; 
              output Core19_Req ; 
              output Core20_Req ; 
              output Core21_Req ; 
              output Core22_Req ; 
              output Core23_Req ; 
              output Core24_Req ; 
              output Core25_Req ; 
              output Core26_Req ; 
              output Core27_Req ; 
              output Core28_Req ; 
              output Core29_Req ; 
              output Core30_Req ; 
              output Core31_Req ; 
              
              output Core0_Addr ;
              output Core1_Addr ;
              output Core2_Addr ;
              output Core3_Addr ;
              output Core4_Addr ;
              output Core5_Addr ;
              output Core6_Addr ;
              output Core7_Addr ;
              output Core8_Addr ;
              output Core9_Addr ;
              output Core10_Addr ; 
              output Core11_Addr ; 
              output Core12_Addr ; 
              output Core13_Addr ; 
              output Core14_Addr ; 
              output Core15_Addr ; 
              output Core16_Addr ; 
              output Core17_Addr ; 
              output Core18_Addr ; 
              output Core19_Addr ; 
              output Core20_Addr ; 
              output Core21_Addr ; 
              output Core22_Addr ; 
              output Core23_Addr ; 
              output Core24_Addr ; 
              output Core25_Addr ; 
              output Core26_Addr ; 
              output Core27_Addr ; 
              output Core28_Addr ; 
              output Core29_Addr ; 
              output Core30_Addr ; 
              output Core31_Addr ; 
              
              
              input Core0_Ack ;
              input Core1_Ack ;
              input Core2_Ack ;
              input Core3_Ack ;
              input Core4_Ack ;
              input Core5_Ack ;
              input Core6_Ack ;
              input Core7_Ack ;
              input Core8_Ack ;
              input Core9_Ack ;
              input Core10_Ack ;
              input Core11_Ack ;
              input Core12_Ack ;
              input Core13_Ack ;
              input Core14_Ack ;
              input Core15_Ack ;
              input Core16_Ack ;
              input Core17_Ack ;
              input Core18_Ack ;
              input Core19_Ack ;
              input Core20_Ack ;
              input Core21_Ack ;
              input Core22_Ack ;
              input Core23_Ack ;
              input Core24_Ack ;
              input Core25_Ack ;
              input Core26_Ack ;
              input Core27_Ack ;
              input Core28_Ack ;
              input Core29_Ack ;
              input Core30_Ack ;
              input Core31_Ack ;
              input  Core0_Data ;
              input  Core1_Data ; 		
              input  Core2_Data ; 
              input  Core3_Data ;
              input  Core4_Data ;
              input  Core5_Data ;
              input  Core6_Data ;
              input  Core7_Data ;
              input  Core8_Data ;
              input  Core9_Data ;
              input  Core10_Data ;
              input  Core11_Data ;
              input  Core12_Data ;
              input  Core13_Data ;
              input  Core14_Data ;
              input  Core15_Data ;
              input  Core16_Data ;
              input  Core17_Data ;
              input  Core18_Data ;
              input  Core19_Data ;
              input  Core20_Data ;
              input  Core21_Data ;
              input  Core22_Data ;
              input  Core23_Data ;
              input  Core24_Data ;
              input  Core25_Data ;
              input  Core26_Data ;
              input  Core27_Data ;
              input  Core28_Data ;
              input  Core29_Data ;
              input  Core30_Data ;
              input  Core31_Data ;

		endclocking
endinterface
