parameter MAX_TEST_COUNT = 5 ;
parameter TEST_COUNT = 2 ;
parameter WAIT_DELAY = 10 ;
`define INTERCONNECT_SINGLE_REQUEST_TEST
`define INTERCONNECT_SINGLE_BANK_MULTIPLE_REQUEST_TEST
